library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity LCL_Project1_14041 is
	
end LCL_Project1_14041;

architecture RTL of LCL_Project1_14041 is
	
begin

	
	
end RTL;
