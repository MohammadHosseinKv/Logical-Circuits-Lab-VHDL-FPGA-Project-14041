LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;


ENTITY LCL_Project1_14041_TB IS
END LCL_Project1_14041_TB;
 
ARCHITECTURE behavior OF LCL_Project1_14041_TB IS 
 
 
    COMPONENT LCL_Project1_14041
    
    END COMPONENT;
    
BEGIN
 
   stim_proc: process
   begin		


      wait;
   end process;

END;
